module cross_correlation (
  input   logic  clk,
  input   logic  reset,

  input   logic  sig_x_i,
  input   logic  sig_y_i,

  output  logic  z_o
);

  // Write your logic here...
  :)

endmodule
